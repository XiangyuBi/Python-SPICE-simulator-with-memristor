

v1 1 0  sin(0 10 20meg)
x1 1 0 1k 16k 14k




.TRAN 0.5n 500n
.Print tran v(1)   i(x1)
.end



